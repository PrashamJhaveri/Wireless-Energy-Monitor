library verilog;
use verilog.vl_types.all;
entity VHDL_vlg_vec_tst is
end VHDL_vlg_vec_tst;
